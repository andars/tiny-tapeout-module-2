localparam PC_FROM_REG   = 2'b00;
localparam PC_FROM_DATA  = 2'b01;

localparam PC_STACK_NOP  = 2'b00;
localparam PC_STACK_PUSH = 2'b01;
localparam PC_STACK_POP  = 2'b10;
